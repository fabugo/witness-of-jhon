module cc(Z, C, S, O, E, C_RE, ZCSO);

	input reg Z, C, S, O, E; // Flag Zero | Flag Carry | Flag Sinal | Flag Overflow | Enable Geral
	input [4:0] C_RE; // Controle RE - Enable Espec�fico: [Z][C][N][O]
	output reg [3:0] ZCSO; // Sa�da das flags

always @(C_RE or E)
	begin
		if(E) 
			case(C_RE)
			 
				5'b01000, 5'b01001: begin // Flag's atualizadas: S, C, Z
					ZCSO[0] = Z;
					ZCSO[1] = C;
					ZCSO[2] = S;					
					end
				
				5'b10001, 5'b10010: begin // Flag's atualizadas: Z, S
					ZCSO[0] = Z;
					ZCSO[2] = S;	
					end
				
				5'b00000, 5'b00001,
				5'b00011, 5'b00100,
				5'b00101, 5'b00110: begin // Flag's atualizadas: Todas
					ZCSO[0] = Z;
					ZCSO[1] = C;
					ZCSO[2] = S;	
					ZCSO[3] = O;	
					end
				
				5'b10001, 5'b10010, 
				5'b10100, 5'b10101, 
				5'b10110, 5'b10111, 
				5'b11000, 5'b11001, 
				5'b11010, 5'b11011, 
				5'b11100, 5'b11101, 
				5'b11110: begin // Flag's atualizadas: Z, S
					ZCSO[0] = Z;	
					ZCSO[2] = S;	
				end
				
				default: begin end // Flag's atualizadas: Nenhuma
			endcase
	end
	
  // * Existe a necessidade do clock?
  // * A justificativa para o uso do enable geral, seria pelo motivo de a atribui��o do estado poder est� sendo feita antes da opera��o ser 
  //   realizada na ULA. Nesse caso, quando a ula finalizar sua opera��o ela poder� mandar um sinal para o RE, habilitando o RE para escrita.
endmodule 