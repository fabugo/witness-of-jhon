// +UEFSHDR----------------------------------------------------------------------
// 2014 UEFS Universidade Estadual de Feira de Santana
// TEC499-Sistemas Digitais
// ------------------------------------------------------------------------------
// TEAM: <Team identification>
// ------------------------------------------------------------------------------
// PROJECT: <Process>
// ------------------------------------------------------------------------------
// FILE NAME  : {module_name}
// KEYWORDS 	: {keywords}
// -----------------------------------------------------------------------------
// PURPOSE: {description}
// -----------------------------------------------------------------------------
// REUSE ISSUES
//   Reset Strategy      : <asychronous, active in low level reset>
//   Clock Domains       : <clock_driver>
//   Instantiations      : <modules_id>
//   Synthesizable (y/n) : <y/n>
// -UEFSHDR----------------------------------------------------------------------
