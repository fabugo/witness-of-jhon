/*
add wave -position insertpoint  \
sim:/IntegracaoModulos/clock
add wave -position insertpoint  \
sim:/IntegracaoModulos/Controle/instrucao
add wave -position insertpoint  \
sim:/IntegracaoModulos/IF/PC/pc_out
add wave -position insertpoint  \
sim:/IntegracaoModulos/ID_RF/A \
sim:/IntegracaoModulos/ID_RF/B \
sim:/IntegracaoModulos/ID_RF/constanteExtendida
add wave -position insertpoint  \
sim:/IntegracaoModulos/EX_MEN/Saida_ULA \
sim:/IntegracaoModulos/EX_MEN/Saida_MemoriaDados
add wave -position insertpoint  \
sim:/IntegracaoModulos/ID_RF/Banco_Registro/registro
add wave -position insertpoint  \
sim:/IntegracaoModulos/EX_MEN/Memoria_Dados/dado_mem
# (vsim-4077) Logging very large object: /IntegracaoModulos/EX_MEN/Memoria_Dados/dado_mem 
*/