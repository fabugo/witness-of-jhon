/*
* @author Patricia Gomes
* @author Kelvin Carmo
* Module: Banco_Registro
* Purpose: Modulo respons�vel por armazenar os registros.
*/

module Banco_Registro (
  Hab_Escrita, // Habilita a escrita no registrador
  Sel_E_SA,    // Endereco da entrada de dados e da saida de dados A, sua fun��o depende do estado de "Hab_Escrita"
  Sel_SB,      // Endereco da saida de dados B
  reset,       // Limpa todos os registros
  clock,       // Pulso de clock
  A,           // Saida A do Banco de Registros
  B,           // Saida B do Banco de Registros
  E);          // Entrada E do Banco de Registros - novo registro a ser armazenado

  parameter bits_palavra = 16;
  parameter end_registros = 3; // Quantidade de bits necess�rios para endere�ar os registros
  parameter num_registros = 8; // Quantidade de registros do Banco de Registros (num_registros = (end_registros^2)-1;)

  output reg [bits_palavra-1:0] A, B;
  input [bits_palavra-1:0] E;

  input [end_registros-1:0] Sel_E_SA, Sel_SB;
  input reset, clock;
  input reg Hab_Escrita;
  reg [bits_palavra-1:0] registro [num_registros-1:0];	// Um vetor de "end_registros" palavras de "bits_palavra" bits

	initial // Inicializa os registradores. // Remover
			begin
			  registro[0] = 16'b0110101111010101;
				registro[1] = 16'b0001110111010110;
				registro[2] = 16'b0001010101101011;
				registro[3] = 16'b0010101011011101;
				registro[4] = 16'b0000000000001101;
				registro[5] = 16'b0000000010101100;
				registro[6] = 16'b0000000000000101;
				registro[7] = 16'b0000000010101011;
<<<<<<< HEAD:rtl/Banco_Registro.sv
			end



	always @(negedge clock, posedge reset) begin

			if(reset) begin
				registro[0] = 16'b0000000000000000;
				registro[1] = 16'b0000000000000000;
				registro[2] = 16'b0000000000000000;
				registro[3] = 16'b0000000000000000;
				registro[4] = 16'b0000000000000000;
				registro[5] = 16'b0000000000000000;
				registro[6] = 16'b0000000000000000;
				registro[7] = 16'b0000000000000000;
			end
			else if(Hab_Escrita) begin
				registro[Sel_E_SA] <= E;
		    end else begin
				A = registro[Sel_E_SA];
				B = registro[Sel_SB];
			end

=======
				registro[8] = 16'b0000000000111111;
				registro[9] = 16'b0001010101100111;
				registro[10] = 16'b0010101010110110;
				registro[11] = 16'b0001110110101111;
				registro[12] = 16'b0000101010000010;
				registro[13] = 16'b0000001101010110;
				registro[14] = 16'b0000110100100111;
				registro[15] = 16'b0011100000100100;
			end

	always_comb
	begin
		//if(!Hab_Escrita)             	// Se a escrita n�o estiver habilitada
			A = registro[Sel_E_SA]; 	// Coloca na sa�da o dado do registrador informado pela entrada Sel_E_SA
		B = registro[Sel_SB]; 			// Coloca na sa�da o dado do registrador informado pela entrada Sel_SB
>>>>>>> origin/mic_arq2:rtl/Banco_Registro.sv
	end

endmodule
