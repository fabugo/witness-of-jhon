
so�ifslkfjsd