/*
*@author Patricia Gomes
*@author Kelvin Carmo
*Module: registers_file
*/
	
module registers_bank #(parameter size_reg=16, addr_reg=2)(/* size_reg = tamanho do dado ( tamanho do registrador) addr_reg = tamanho do endere�o do registrador*/
	input [addr_reg-1:0] addr_A, //endere�o do registrador onde o operando A ser� gravado.
	input [addr_reg-1:0] addr_B, //endere�o do registrador onde o operando B ser� gravado.
	input [addr_reg-1:0] addr_R,//endere�o do registrador onde o dado ser� gravado.
	input write_reg, //habilitador de escrita.
	input clock,
	input reset,
	input [size_reg-1:0] write_data, //dado.
	output reg [size_reg-1:0] data_A, //dado que sai do registrador A.
	output reg [size_reg-1:0] data_B); //dado que sai do registrador B.

	reg [size_reg-1:0] registers[0:(1'b1 << addr_reg)-1];//2^N registradores de M bits
			
	initial // innicializa os registradores.
			begin
				registers[0] = 16'b0000000000000000;
				registers[1] = 16'b0000000000000000;
				registers[2] = 16'b0000000000000000;
				registers[3] = 16'b0000000000000000;
			end

	always_comb 
		begin
			data_A = registers[addr_A]; //coloca na sa�da o dado do registrador informado pela entrada addr_A
			data_B = registers[addr_B]; //coloca na sa�da o dado do registrador informado pela entrada addr_B
		end

	always@(posedge clock, negedge reset) 
		begin// sinal de escrita ou leitura
			if(!reset) //Reset ass�ncrono
				begin 
					registers[0] = 16'b0000000000000000;
					registers[1] = 16'b0000000000000000;
					registers[2] = 16'b0000000000000000;
					registers[3] = 16'b0000000000000000;
				end
			else if(write_reg) 
				registers[addr_R] <= write_data;//*escreve o dado no registrador destino, de endere�o informado pela entrada "addr_R"
		end
	 
endmodule